library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

entity ramBlock is
port (clk :in std_logic;
	addr: in std_logic_Vector(12 downto 0);
	output : out std_logic_vector(7 downto 0));
	
end ramBlock;

architecture Behavioral of ramBlock is
type arr is array (0 to 7999) of integer range 0 to 255;
constant data8KB:arr:=(127, 127, 126, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 127, 127, 126, 127, 126, 126, 126, 125, 125, 125, 125, 125, 125, 125, 125, 125, 124, 124, 124, 124, 124, 124, 125, 124, 124, 124, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 125, 125, 125, 125, 126, 126, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 122, 122, 122, 122, 122, 122, 122, 122, 121, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 121, 121, 121, 121, 121, 121, 121, 122, 122, 122, 121, 121, 121, 121, 121, 121, 121, 121, 122, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 120, 121, 121, 121, 121, 121, 121, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 121, 121, 120, 120, 120, 121, 121, 121, 120, 120, 120, 120, 120, 120, 120, 120, 121, 121, 120, 121, 121, 121, 121, 121, 121, 121, 121, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 121, 121, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 121, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 126, 126, 125, 126, 126, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 126, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 127, 127, 128, 127, 127, 127, 127, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 127, 127, 127, 127, 128, 128, 128, 128, 128, 127, 127, 127, 127, 127, 128, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 127, 127, 128, 128, 127, 127, 127, 128, 128, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 127, 128, 128, 128, 127, 127, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 127, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127,
127, 128, 128, 128, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 127, 127, 127, 127, 127, 126, 126, 126, 126, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 127, 127, 128, 129, 129, 130, 131, 132, 132, 133, 134, 135, 136, 136, 137, 138, 138, 138, 138, 139, 138, 138, 137, 136, 135, 133, 131, 130, 128, 126, 124, 123, 121, 120, 119, 118, 117, 116, 116, 116, 116, 116, 117, 117, 118, 118, 119, 120, 120, 120, 121, 121, 121, 122, 122, 123, 123, 123, 124, 125, 126, 127, 128, 129, 131, 132, 134, 136, 138, 139, 141, 142, 143, 145, 145, 145, 145, 145, 144, 143, 141, 138, 135, 134, 132, 128, 127, 127, 123, 121, 121, 119, 117, 118, 119, 118, 119, 120, 119, 119, 120, 119, 119, 120, 119, 118, 118, 117, 115, 115, 117, 116, 116, 118, 119, 119, 121, 122, 122, 125, 126, 127, 129, 130, 130, 131, 133, 134, 136, 138, 139, 141, 143, 145, 146, 149, 151, 152, 153, 152, 150, 145, 141, 139, 137, 133, 132, 133, 129, 124, 122, 120, 115, 115, 117, 117, 119, 122, 122, 122, 123, 123, 122, 122, 121, 120, 120, 118, 116, 116, 116, 115, 116, 118, 116, 116, 118, 118, 118, 122, 124, 124, 126, 128, 128, 128, 130, 130, 132, 135, 136, 138, 141, 143, 144, 148, 150, 152, 156, 157, 157, 156, 149, 142, 142, 140, 130, 130, 136, 129, 122, 124, 120, 111, 114, 118, 115, 117, 124, 123, 122, 127, 125, 123, 126, 124, 118, 118, 118, 112, 110, 113, 110, 108, 111, 110, 108, 110, 111, 110, 114, 118, 118, 120, 124, 124, 124, 127, 128, 129, 134, 136, 136, 140, 143, 143, 145, 150, 151, 153, 158, 160, 160, 162, 160, 149, 145, 146, 139, 129, 133, 136, 128, 125, 127, 119, 111, 116, 116, 113, 118, 124, 122, 123, 126, 123, 122, 125, 121, 117, 118, 115, 108, 107, 109, 104, 104, 106, 104, 104, 106, 105, 106, 112, 114, 115, 120, 123, 122, 124, 127, 126, 129, 134, 135, 137, 142, 144, 144, 147, 150, 152, 156, 160, 161, 163, 165, 166, 163, 154, 148, 146, 138, 130, 131, 134, 128, 125, 127, 119, 111, 114, 116, 114, 118, 125, 126, 127, 131, 128, 125, 127, 124, 120, 119, 113, 106, 104, 103, 97, 99, 103, 101, 101, 105, 104, 104, 110, 113, 114, 120, 124, 122, 124, 127, 127, 129, 135, 137, 138, 143, 143, 143, 146, 149, 150, 154, 158, 159, 162, 165, 165, 167, 170, 159, 151, 150, 140, 126, 125, 128, 123, 119, 124, 118, 108, 109, 109, 108, 113, 121, 125, 128, 133, 131, 129, 132, 128, 124, 123, 118, 110, 104, 99, 92, 90, 92, 90, 93, 100, 100, 101, 107, 112, 116, 124, 130, 131, 134, 135, 132, 132, 135, 136, 138, 143, 143, 142, 144, 144, 144, 147, 152, 154, 157, 162, 163, 165, 169, 170, 171, 164, 153, 147, 136, 123, 115, 118, 119, 115, 117, 115, 105, 103, 103, 104, 110, 121, 132, 137, 143, 143, 138, 138, 131, 126, 123, 117, 110, 100, 95, 87, 82, 85, 84, 88, 96, 101, 106, 112, 121, 126, 132, 140, 141, 142, 142, 139, 137, 136, 136, 137, 139, 141, 140, 140, 140, 140, 143, 147, 150, 154, 159, 161, 163, 167, 169, 170, 176, 167, 151, 143, 128, 108, 103, 103, 105, 109, 115, 117, 108, 108, 107, 107, 121, 129, 142, 152, 155, 151, 140, 133, 118, 107, 105, 93, 86, 83, 75, 72, 73, 81, 87, 99, 115, 120, 129, 137, 137, 140, 141, 140, 134, 131, 124, 113, 111, 109, 109, 119, 128, 136, 143, 150, 152, 152, 158, 158, 160, 164, 163, 159, 157, 155, 151, 152, 155, 159, 156, 139, 130, 115, 93, 93, 98, 110, 129, 138, 146, 135, 128, 122, 111, 126, 131, 142, 154, 149, 140, 121, 108, 93, 81, 89, 85, 87, 97, 93, 97, 104, 114, 123, 134, 145, 142, 136, 133, 120, 115, 116, 113, 111, 111, 107, 99, 103, 110, 118, 135, 152, 161, 166, 166, 158, 150, 147, 141, 138, 140, 138, 135, 137, 140, 143, 155, 169, 178, 188, 199, 172, 141, 130, 88, 63, 81, 89, 114, 148, 159, 153, 135, 132, 107, 108, 137, 133, 151, 160, 142, 118, 103, 94, 75, 88, 110, 96, 110, 113, 94, 101, 114, 125, 128, 144, 143, 117, 112, 105, 87, 103, 115, 111, 111, 112, 96, 90, 112, 126, 141, 172, 176, 163, 157, 137, 116, 112, 121, 120, 131, 150, 150, 151, 166, 164, 160, 171, 177, 170, 178, 193, 161, 123, 122, 73, 41, 79, 91, 122, 178, 189, 174, 148, 137, 96, 87, 135, 124, 146, 168, 142, 114, 103, 97, 77, 97, 127, 99, 107, 105, 69, 79, 108, 129, 147, 177, 168, 125, 107, 83, 54, 76, 102, 106, 121, 134, 113, 111, 136, 143, 153, 176, 164, 134, 122, 103, 89, 106, 134, 146, 164, 175, 159, 145, 151, 145, 147, 162, 171, 171, 177, 181, 189, 168, 120, 115, 69, 33, 72, 96, 139, 205, 217, 197, 152, 122, 77, 56, 116, 112, 142, 170, 145, 119, 105, 104, 86, 102, 130, 87, 86, 87, 56, 87, 134, 165, 183, 199, 158, 95, 62, 30, 23, 69, 116, 143, 163, 169, 134, 119, 127, 112, 124, 133, 123, 110, 112, 113, 116, 144, 156, 154, 163, 145, 128, 124, 129, 137, 154, 176, 179, 186, 191, 178, 191, 180, 99, 100, 77, 17, 72, 124, 152, 225, 243, 194, 126, 90, 56, 24, 122, 141, 153, 197, 164, 119, 104, 111, 89, 95, 136, 78, 57, 79, 54, 93, 169, 205, 198, 201, 142, 46, 22, 10, 14, 88, 157, 178, 189, 188, 130, 88, 100, 78, 88, 120, 120, 117, 135, 140, 131, 151, 154, 130, 135, 127, 113, 123, 139, 152, 168, 190, 185, 179, 178, 168, 160, 182, 182, 107, 102, 99, 18, 72, 139, 149, 231, 248, 181, 114, 73, 53, 33, 140, 173, 162, 203, 152, 108, 95, 110, 104, 102, 136, 74, 41, 74, 62, 114, 196, 221, 196, 176, 104, 15, 15, 21, 52, 134, 185, 190, 178, 153, 96, 58, 76, 66, 90, 127, 129, 134, 146, 142, 124, 135, 131, 110, 128, 130, 126, 146, 155, 156, 169, 181, 159, 164, 169, 156, 160, 178, 194, 131, 97, 114, 37, 59, 150, 150, 212, 243, 173, 107, 70, 62, 47, 132, 189, 150, 186, 151, 107, 105, 123, 120, 98, 117, 66, 21, 72, 88, 133, 209, 228, 179, 140, 94, 5, 12, 50, 69, 131, 188, 179, 155, 142, 93, 46, 65, 73, 83, 132, 150, 141, 149, 147, 115, 119, 128, 117, 132, 148, 141, 146, 151, 155, 167, 179, 175, 171, 166, 163, 164, 185, 216, 147, 108, 118, 33, 45, 142, 158, 213, 254, 176, 95, 59, 54, 47, 140, 200, 158, 185, 149, 107, 109, 131, 126, 96, 106, 55, 19, 80, 109, 155, 218, 218, 153, 111, 71, 13, 26, 61, 94, 133, 177, 178, 152, 143, 95, 46, 51, 59, 90, 135, 170, 162, 151, 138, 102, 108, 122, 131, 148, 154, 150, 144, 146, 152, 163, 177, 173, 172, 160, 169, 171, 193, 210, 107, 80, 85, 14, 79, 175, 191, 234, 230, 131, 50, 43, 60, 71, 183, 194, 149, 168, 135, 116, 128, 150, 106, 64, 65, 13, 29, 119, 157, 192, 225, 180, 95, 79, 49, 30, 69, 81, 96, 136, 164, 159, 158, 144, 88, 49, 46, 50, 94, 151, 171, 165, 154, 122, 101, 118, 124, 130, 143, 135, 132, 143, 155, 162, 169, 171, 156, 157, 160, 164, 175, 196, 209, 125, 58, 87, 50, 76, 183, 194, 208, 217, 135, 64, 49, 79, 84, 156, 197, 144, 156, 146, 133, 129, 142, 109, 50, 61, 45, 55, 134, 175, 182, 191, 168, 91, 71, 74, 49, 71, 103, 116, 132, 167, 162, 133, 123, 83, 45, 60, 90, 111, 144, 158, 133, 127, 130, 118, 129, 140, 129, 126, 131, 132, 147, 167, 172, 170, 168, 158, 143, 150, 168, 174, 182, 205, 207, 106, 73, 99, 44, 99, 195, 186, 216, 208, 115, 52, 56, 85, 94, 189, 189, 142, 160, 147, 127, 127, 138, 81, 48, 70, 53, 85, 153, 167, 152, 164, 130, 68, 88, 83, 58, 81, 109, 103, 129, 171, 141, 119, 107, 58, 41, 77, 104, 116, 150, 143, 116, 131, 131, 120, 133, 137, 118, 126, 144, 148, 154, 167, 163, 154, 158, 157, 148, 154, 167, 168, 183, 214, 187, 93, 95, 86, 53, 136, 188, 185, 212, 167, 89, 54, 80, 101, 135, 199, 155, 138, 146, 137, 127, 130, 117, 60, 59, 72, 75, 118, 155, 146, 135, 143, 105, 90, 103, 89, 78, 81, 103, 113, 138, 156, 132, 109, 90, 64, 60, 88, 107, 116, 133, 132, 125, 137, 139, 128, 130, 127, 122, 133, 146, 156, 155, 158, 157, 148, 151, 167, 163, 166, 181, 178, 184, 213, 194, 88, 87, 107, 76, 129, 183, 173, 186, 171, 98, 62, 89, 106, 121, 183, 154, 125, 149, 153, 134, 132, 118, 57, 54, 81, 87, 113, 145, 130, 118, 139, 118, 95, 106, 91, 70, 78, 102, 115, 139, 152, 127, 105, 94, 68, 59, 85, 99, 114, 133, 136, 132, 143, 139, 127, 130, 127, 127, 139, 151, 159, 160, 153, 149, 159, 163, 167, 170, 164, 164, 180, 187, 196, 181, 96, 89, 118, 101, 125, 168, 166, 168, 148, 111, 76, 98, 117, 121, 152, 135, 125, 143, 163, 143, 120, 105, 67, 62, 91, 101, 102, 122, 118, 116, 141, 133, 110, 107, 99, 84, 83, 93, 112, 133, 137, 126, 112, 103, 86, 72, 80, 91, 108, 128, 139, 141, 143, 142, 137, 138, 134, 132, 135, 139, 147, 152, 151, 156, 166, 161, 162, 166, 160, 157, 174, 182, 196, 182, 105, 96, 124, 117, 122, 149, 149, 147, 138, 122, 98, 109, 119, 118, 139, 130, 125, 139, 160, 142, 122, 116, 94, 87, 100, 99, 91, 106, 111, 119, 143, 141, 119, 111, 108, 99, 92, 93, 99, 115, 122, 116, 112, 118, 106, 91, 88, 90, 98, 114, 125, 125, 131, 135, 137, 143, 139, 131, 127, 128, 132, 138, 151, 155, 159, 161, 163, 161, 157, 149, 154, 170, 176, 186, 169, 123, 121, 142, 123, 111, 125, 129, 141, 140, 127, 108, 119, 127, 131, 141, 129, 116, 127, 140, 132, 133, 131, 115, 104, 110, 100, 92, 96, 99, 107, 125, 129, 123, 126, 122, 115, 106, 95, 91, 106, 113, 105, 106, 114, 111, 101, 100, 97, 100, 108, 109, 109, 115, 125, 136, 147, 147, 138, 132, 130, 128, 133, 139, 143, 146, 145, 148, 153, 157, 152, 150, 154, 160, 168, 178, 183, 177, 164, 154, 146, 133, 125, 134, 140, 127, 121, 122, 121, 127, 135, 127, 114, 114, 115, 124, 135, 132, 127, 126, 121, 119, 122, 117, 106, 103, 107, 108, 111, 113, 111, 109, 110, 108, 104, 104, 105, 102, 100, 101, 101, 100, 100, 100, 98, 99, 101,
104, 109, 114, 118, 121, 123, 125, 131, 137, 141, 145, 147, 147, 148, 153, 156, 156, 155, 155, 154, 157, 164, 169, 171, 174, 175, 172, 164, 153, 154, 162, 155, 138, 140, 142, 133, 132, 126, 113, 109, 112, 112, 113, 113, 109, 112, 117, 117, 117, 122, 123, 120, 120, 116, 110, 108, 110, 110, 106, 103, 100, 99, 101, 100, 96, 99, 101, 99, 101, 104, 103, 102, 104, 107, 109, 112, 113, 112, 113, 116, 121, 129, 132, 135, 139, 140, 142, 145, 147, 150, 152, 154, 155, 157, 159, 161, 164, 165, 163, 157, 157, 164, 171, 171, 162, 153, 156, 161, 150, 138, 137, 131, 124, 120, 115, 111, 114, 114, 110, 107, 104, 105, 112, 114, 113, 114, 115, 116, 118, 117, 113, 108, 106, 105, 104, 104, 102, 101, 102, 105, 103, 100, 105, 111, 110, 107, 109, 112, 112, 114, 115, 115, 116, 116, 118, 121, 125, 129, 133, 133, 133, 135, 140, 144, 146, 147, 148, 152, 158, 160, 159, 157, 154, 153, 156, 158, 159, 161, 164, 167, 166, 157, 147, 148, 150, 144, 134, 129, 129, 126, 121, 115, 109, 106, 106, 106, 105, 103, 103, 109, 114, 115, 116, 116, 117, 118, 117, 114, 113, 111, 110, 111, 108, 106, 106, 107, 109, 108, 106, 109, 110, 109, 112, 114, 112, 112, 114, 114, 116, 118, 118, 119, 120, 122, 125, 127, 128, 130, 134, 138, 141, 144, 146, 148, 149, 150, 150, 149, 148, 149, 152, 155, 154, 151, 151, 154, 155, 153, 152, 154, 152, 145, 141, 144, 141, 129, 127, 129, 125, 120, 117, 113, 113, 116, 115, 114, 113, 111, 115, 120, 119, 116, 117, 117, 117, 117, 116, 114, 112, 112, 112, 111, 110, 107, 107, 111, 112, 107, 107, 111, 113, 113, 113, 112, 114, 117, 117, 117, 119, 119, 120, 124, 126, 127, 129, 132, 133, 136, 138, 139, 142, 145, 147, 148, 150, 151, 148, 150, 153, 151, 148, 150, 150, 149, 150, 150, 149, 149, 151, 150, 142, 139, 142, 140, 133, 130, 129, 128, 127, 122, 119, 118, 117, 116, 114, 110, 108, 110, 111, 109, 110, 111, 111, 112, 112, 110, 108, 106, 105, 104, 105, 104, 102, 103, 107, 107, 104, 105, 107, 109, 111, 112, 113, 115, 118, 121, 124, 126, 127, 128, 130, 132, 134, 137, 139, 141, 143, 143, 144, 147, 150, 151, 151, 151, 151, 152, 152, 151, 151, 150, 149, 149, 148, 148, 149, 148, 148, 146, 141, 140, 141, 139, 134, 132, 131, 128, 126, 122, 118, 116, 114, 112, 111, 108, 107, 109, 112, 112, 111, 110, 110, 109, 110, 108, 107, 107, 108, 108, 107, 106, 105, 104, 106, 107, 106, 109, 112, 114, 116, 119, 120, 124, 127, 128, 129, 130, 131, 134, 136, 137, 137, 138, 139, 140, 142, 143, 144, 144, 145, 145, 146, 147, 148, 147, 145, 144, 144, 144, 143, 141, 140, 139, 139, 139, 138, 139, 139, 137, 135, 135, 136, 134, 130, 126, 126, 125, 122, 120, 121, 120, 118, 117, 115, 112, 109, 108, 108, 109, 110, 109, 109, 109, 109, 108, 107, 106, 108, 109, 109, 109, 109, 111, 113, 114, 115, 116, 118, 120, 121, 122, 124, 126, 128, 128, 129, 129, 131, 132, 133, 134, 134, 134, 135, 136, 137, 137, 138, 139, 139, 140, 140, 140, 141, 142, 141, 140, 139, 139, 139, 139, 139, 137, 137, 137, 137, 137, 136, 135, 135, 135, 135, 135, 135, 134, 132, 131, 130, 128, 126, 126, 124, 123, 123, 122, 118, 116, 116, 115, 114, 114, 113, 112, 113, 114, 113, 113, 113, 112, 112, 112, 113, 114, 116, 117, 119, 120, 121, 121, 122, 122, 123, 124, 124, 123, 124, 126, 127, 128, 130, 130, 130, 130, 130, 131, 133, 133, 133, 133, 134, 135, 134, 135, 136, 136, 136, 136, 135, 135, 135, 135, 135, 136, 136, 138, 139, 138, 136, 137, 136, 134, 135, 135, 133, 134, 134, 133, 133, 134, 132, 129, 127, 125, 124, 123, 122, 121, 121, 120, 119, 118, 117, 116, 114, 113, 113, 113, 114, 116, 116, 115, 116, 116, 116, 117, 117, 117, 117, 118, 119, 120, 121, 122, 121, 122, 122, 122, 123, 124, 125, 126, 127, 127, 127, 127, 128, 128, 129, 130, 130, 130, 131, 131, 131, 131, 133, 134, 134, 135, 136, 136, 137, 138, 138, 138, 138, 138, 138, 138, 139, 139, 138, 137, 136, 134, 132, 131, 131, 131, 130, 129, 128, 128, 127, 126, 125, 123, 122, 122, 122, 121, 121, 122, 122, 121, 120, 119, 118, 119, 119, 117, 117, 118, 118, 118, 118, 117, 116, 117, 116, 116, 116, 117, 118, 118, 118, 118, 118, 120, 121, 122, 122, 124, 125, 126, 127, 128, 129, 129, 130, 130, 131, 131, 132, 133, 135, 135, 135, 136, 136, 137, 137, 137, 138, 139, 140, 139, 138, 137, 137, 137, 137, 136, 135, 134, 133, 133, 132, 131, 130, 130, 128, 127, 126, 126, 126, 126, 125, 124, 123, 122, 121, 121, 121, 120, 120, 121, 121, 120, 119, 119, 119, 118, 117, 117, 118, 118, 118, 118, 118, 118, 118, 118, 117, 117, 118, 120, 121, 122, 123, 123, 123, 124, 125, 126, 127, 129, 130, 130, 131, 132, 133, 133, 133, 133, 134, 135, 135, 136, 136, 136, 136, 135, 135, 135, 136, 135, 135, 135, 134, 133, 133, 133, 132, 131, 130, 129, 129, 129, 129, 128, 128, 128, 126, 125, 124, 124, 125, 124, 124, 124, 123, 122, 122, 122, 121, 121, 121, 120, 120, 119, 119, 119, 120, 120, 120, 119, 118, 118, 119, 119, 119, 120, 121, 122, 122, 123, 124, 124, 125, 126, 127, 127, 128, 129, 130, 130, 130, 131, 131, 132, 133, 133, 133, 133, 134, 134, 134, 135, 135, 134, 134, 134, 134, 134, 134, 134, 134, 133, 132, 132, 131, 131, 131, 131, 130, 129, 129, 128, 128, 127, 127, 126, 126, 125, 124, 124, 124, 123, 123, 123, 122, 121, 120, 120, 120, 120, 120, 120, 118, 118, 118, 119, 118, 118, 119, 119, 119, 119, 119, 119, 120, 122, 122, 123, 123, 123, 124, 125, 126, 126, 126, 127, 128, 128, 129, 130, 130, 131, 131, 132, 132, 132, 132, 133, 133, 133, 134, 134, 134, 134, 134, 133, 133, 133, 132, 132, 132, 131, 131, 130, 129, 129, 129, 128, 127, 126, 126, 126, 125, 125, 125, 124, 124, 123, 122, 121, 122, 122, 122, 122, 122, 121, 121, 121, 120, 120, 120, 120, 121, 121, 120, 121, 121, 121, 121, 122, 122, 123, 124, 124, 125, 126, 126, 127, 128, 128, 128, 129, 130, 130, 131, 131, 131, 131, 132, 132, 133, 133, 133, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 133, 133, 133, 132, 132, 131, 130, 130, 129, 129, 129, 128, 127, 127, 126, 126, 125, 125, 124, 123, 122, 122, 122, 122, 121, 121, 120, 120, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 120, 120, 120, 120, 121, 121, 122, 123, 124, 124, 124, 124, 125, 126, 126, 127, 128, 128, 128, 129, 129, 129, 130, 131, 131, 131, 132, 132, 132, 132, 132, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 132, 132, 131, 131, 130, 130, 129, 128, 128, 127, 127, 126, 126, 125, 125, 124, 124, 124, 123, 123, 123, 122, 122, 122, 122, 122, 121, 121, 121, 121, 121, 121, 122, 121, 121, 121, 121, 120, 121, 122, 122, 123, 123, 123, 123, 124, 125, 126, 126, 127, 127, 127, 128, 129, 130, 131, 131, 132, 132, 132, 132, 133, 133, 133, 134, 134, 134, 134, 134, 134, 134, 134, 133, 133, 133, 132, 132, 132, 132, 132, 131, 130, 129, 129, 128, 128, 127, 126, 126, 125, 125, 124, 124, 124, 124, 123, 122, 122, 122, 122, 121, 121, 121, 121, 121, 121, 121, 121, 121, 120, 120, 120, 121, 121, 121, 121, 121, 121, 121, 122, 122, 123, 123, 124, 125, 125, 126, 127, 127, 127, 128, 128, 129, 130, 130, 131, 131, 130, 130, 131, 131, 132, 132, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 132, 131, 131, 131, 130, 130, 130, 130, 129, 128, 128, 127, 127, 126, 126, 126, 125, 125, 124, 124, 123, 123, 122, 122, 122, 122, 121, 121, 120, 120, 120, 121, 120, 120, 120, 120, 120, 120, 120, 121, 121, 121, 122, 122, 122, 123, 124, 124, 124, 125, 125, 126, 127, 128, 128, 128, 129, 129, 129, 130, 130, 131, 132, 132, 132, 132, 133, 133, 133, 133, 133, 133, 133, 133, 132, 132, 132, 131, 131, 131, 130, 130, 130, 129, 129, 128, 128, 127, 127, 127, 126, 126, 126, 125, 124, 124, 124, 124, 124, 124, 123, 123, 123, 122, 122, 123, 123, 123, 122, 122, 122, 123, 123, 122, 122, 122, 122, 122, 122, 123, 123, 123, 124, 124, 124, 124, 125, 126, 126, 127, 127, 127, 128, 128, 128, 129, 129, 129, 130, 130, 130, 130, 129, 129, 130, 130, 130, 130, 130, 130, 130, 130, 130, 129, 129, 129, 129, 129, 129, 129, 128, 128, 128, 128, 128, 127, 128, 128, 127, 127, 127, 127, 126, 126, 126, 126, 125, 125, 125, 125, 124, 124, 124, 124, 124, 124, 124, 124, 123, 123, 124, 124, 124, 124, 124, 124, 124, 124, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 128, 128, 129, 128, 128, 128, 128, 128, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 125, 125, 125, 125, 125, 125, 124, 124, 125, 124, 124, 124, 124, 124, 124, 125, 125, 124, 124, 124, 125, 125, 126, 126, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 129, 128, 128, 128, 128, 128, 128, 128, 128, 128, 129, 129, 128, 128, 128, 128, 128, 128, 128, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 125, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 129, 129, 129, 129, 129, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 127, 128, 128, 128, 128, 128, 127, 126, 126, 127, 127, 127, 127, 127, 127, 126, 125, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127,
127, 126, 126, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 126, 127, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 126, 126, 127, 127, 127, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 127, 126, 126, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 127, 127, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 126, 127, 127, 127, 127, 127, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 127, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 126, 127, 126, 126, 126, 127, 127, 127, 126, 126, 126, 127, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 126, 127, 127, 127, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 127, 126, 127, 127, 127, 126, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 126, 127, 127, 127, 127, 126, 126, 127, 126, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 126, 127, 127, 127, 126, 126, 126, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 127, 127, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 127, 126, 126, 126, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 126, 127, 127, 127, 126, 126, 126, 126, 126, 126, 126, 127, 126, 127, 127, 127, 127, 127, 126, 126, 126, 126, 126, 127, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 126);

begin
process(clk)
begin
	-- Data is stored in the above array. Data corresponding to inputted address is sent to top module.
	if(rising_edge(clk)) then
		output <= conv_std_logic_vector(data8KB(conv_integer(addr)),8);
	end if;
end process;
end Behavioral;